BZh91AY&SY�; u߀Rxg����������P��ݩu�7v�ܺw7	DSii����= M  42�JL&H ��=@���@  �ЈM!�=��OD��H� h ��dd2`��&�F�@�&F 	$	��F����ɒz#�=M @h4mLQI3&9�3��p
B��|?{tM!�7�B�fvS;��v��IX��!iF�Z�X���E��T���Jm%��Klh�ͳ+�k���\�7~�z�!�S�w�wstn�v�BYn���*^q)���� �o�3��4T4\]$���"�9e�_ӣ����YZ�Т�����n k�HM��}�r�ಇIR����� �&l`�:��6������zsk�V��^�V,��)i7����x�*�U�I:I-�����a�u}�j�	)���a�[�tI!�sY ���U
.v�LT�{�W0i(��\��wȫJ1��������&8��M�f?9,��0���se߳g[;	�h����������8�FZ����[�U4ι�����ڎ���1�l%�-�]+Z�����`J��ݣ���Zku[BنS�H6�G�xߓ����b鈇z<��s��`>�U�A�d����2�%Q 0в]6����Rx���C33�3�,Yo
ϳn@�H������J�����M5���ȂY�5lg\�X��7؄�H�
Xd�Bʫ�=�%�mS�$���m�㘿��h,9ا�b>��Q�D�r��d��.�"�E+��C2]�@{b��c�ݒ'vݾ�d%�yV֋��
���ПDk����/��E�Wt���x�����)����n�VӘdWb�,�J��I�w� 2�12���̈pL�'���`\����!�@����6���:s*�=G
�0.�N��W�5�I�ى"�73Д�D}^�`A=�l�71�M��{�FAִT��ji�d}�	1w��L �ck�$zF����B�!b�I�~�sp�u��@5��C�鍜>2(�g�yIX,��m����`ɟ^g�
8bDU�:�����F����%�,a�z<�b-�J�ȣ�ʖ,��ueiK��]M�W
�^c��p�EU�pT��Ր�8� ���N���ƟT���]t��^FM��~P�F�C���%c����H�
Ag`