BZh91AY&SY#�~� �߀Rxg����������P޸�7p�if��H�@56�����6P=M�h4���'����mA�  �    %4!
zF�'�MM��'��A�� F���!�	�4ѣ4ɑ� �H���0L��S��z(ɲ�mA��� ��$����:�N!DT$��G���?�+v�����۩����9�uW��:XE�L�~�Zj !�e�
�_W:c��\1G7�V��X�g���6~X��HC�<m����i�ws�9�ܝ6K*�p$�_λ/&�͌K�N��BEU�(�U4H@D� ��������UEg�+Y�^��h+
��{���w�ACA(�Ы鄘�5gs�[v�L߽,E������!�.�x/�S�Ʒ:)(��w���h;G��I��'I%��x���9COk~�
�JiAe�"]��	��B5�R�W�.Yc�����iWbLf���pL!J!	��y��֧M���y�Ť��c���I�%3�R�d�-�����D@��p,-�Jz켶����N1�n��t<k�=枓9i��\�瀽�r�T�}�Bt���|�uCo ј;�B�f!Σg�d��u��fm#�c��5<�)Y�hک�	�}/H�񉧃`p0�Y�rdf�Ry��҆fg�gM,Ǵ�w�^P�9�@=v87�[D�E��iz��yd����쇌'����2�6��E���B	`C��|����;K��ZOM ���6�5�*�>dq���Z�S9�b`�2��B�㌘;�Ec�-��_>��̛x3#��yK֞(��eL�r�2j	� �(#{5Gq�^6�ãǁ�dj����|�&��]R]��eC���ds@ Jwa�L��&L�F��۷�-))8�PQ^���=��X`b�!@�q��g�V�X��8��!�'�H�����%��%��M���mu� �(Z��d����g��k��,8G).s`/�4�6Dhˡj��:6#�
\�֑謴��i�{�-���r&'E�'&9��1�6j RV%˶H(#4�1P2}Y�'x�6E�<�ӯuSy��1�2��7�hن8L`ZT]1rZ�z�j+Fv"[S���zHw|����ќ�c��D����/��m�Qy"D���ɰ��Zb̋!Cj�����7�#��2[���.�p� Gx��