BZh91AY&SYbJ�q ߀Px�׿�߰����P~t����4B���4�4    �DM4�=Q��?Tɐ�z�D�!��`%4�Bi4��F�   4 sFLL LFi�#ɀF	"M2M2hL�4�=54�@hF@cQ��m(��J@:C�^(2��d'dv�pT�K{F,`�Z��A��I������q*dd����h�Tg�*ɥPʺJ�Y�E�!*lpAa:n�5WVI�^mG��Q1��(a0�yY�s吇L���	���$�CfDA`S\��Yp��-�٨�O�`B*�C�����6�I}a����=���,�H��2�-�taCV��%�"<T"af&1O=��r�\��!#�>����M��F����qA6�h6�	�
K� މ!�@us	��YI���3!Q�r��.�~NP�j�`�;F�$'�)�N�*"�,�#|�2LmǓH����ɜ[qT	���CQ�\i+yc��uj]�=���ý��	��rWc�U�k����%``'
T`GtHT�W�A��*F;��7"���-�A�5��[�\P��D
�K��*V�2y,������,�"���{�#!um\c\�@������FЂ1�{FL8�plT�br���$ ��z��8�,@�&P�)u�0<���h��x�l���x�hd�s�t���zmK�;��v��:Am9��Y40�.c�-! ���5h�30�D��h}::�B�7�M!�!E*PƮp+�9h¼j+qMP�E]��:��~�*3�.�<�q��,2YTcK�kn�Z?��"�(H1%c��