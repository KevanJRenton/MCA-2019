BZh91AY&SY�4��  �_�Pxc����߰����P8��ެ�s����������F�F��4 24&�=@�H�MD�A�     "$4B�&iL�4 OH�L�1�2`� 4a�JoT����Q��L�� Che��B VbT!�����hm�"}{.`u4s�k��\Y��8�䗰�����[q\WI�ץ�ۂ*q�
2��+����rII���^И߻��*�������Yo*#s�VSD�K9H7:<��52Y����N�V�2�4�dվm�/=�5Ǚb�ӵ��3�aȎ�m���[b�ӑ�⤔���;,/r�^3c��$��3t�w2��y��u��멗^U�o�]��^�6h�r��P�q���<uG&ÍՍa�:�F,ܡS�6*"̹Y{��ʳ����L8�ń�F�NV�+Q��Ǩ�3?�^�SlA�	o��#KA�4J��3
����4�������J�t�]9�C��@&qDvd�\Nzl��<8�\�ƁS�0�gZ=��M�]<��,���u�$�h�5�q�i&T���:��S䆂r*x�㴩l�//�:�3*��)��ρ55��b����t��1m�B�guj�Bj��"�Q�H�Ӆ�a�����nE�aE�dw,��Em�o&�W��b���Ğz�d�ʈ:�(���~�p�I9Ϭ���S;Qn4\�*� `*B�$A )BC ma��Eڤ	
@�s2%e�r�m�oF�g����CE���=Q3��.W����3g+�B�.)}��BtIҪ���8�����L.R��aq���"�v��;�BOU�rE8P��4��