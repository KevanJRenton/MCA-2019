BZh91AY&SYA=+8 �߀Ryg����������PޮR�wp��fe�$�)? *~���Ƃ�� �C#�Sj�L�@    � )�	1�i��3���$ښhd��z�q�&�CL	��14�@IB2m$��������@ 4=F��$̆1gф�A%ZIR(�q�Ri������x��ľ1ƪ.�����+��3eAU)0C��l�s���p�0��j;�]���cy�Ѫm��R��O3�jAg����m�K�B7�9]ܷ�MS�bY�͗�R���~a5�K�@�! ]D sn<;�/��ʛ�Mvl��ٰHB��s�����rp6)L�l`��Q��r@�[�k��~��v�D�f�l�>T�w�!�ᣐ�%�޲�4�+&V:�&qz�	#q$�$��'�9_F��7y���T%4� ���w��\&C�=0d�H��L�9=��z��*�]��dF��C,�m�b���if��T,8,�)]ur��_uA��j�tI;"3�����q�47�p�9����L���jg�͚��U�����镟4s<] eD����@6�xn��0ѐ5|��os����$�M�؍m�bt1��^?+i�T�ҿ��P�w�8�KVk9Y����贡����&z�f>��>M+�8[�	�v=}V8�.ꤑP�r���$�yd����쇌�vP��2���r���JGh�0%�'E�g��Bn��ɲ��{0�QX�c�'�F�Z���'<棡	6=�N^���.�6g�7�գag���Ĥ��D�1Z�aB�L��#N���4���c`�l�Q���/�a���28P5��Tw5������p3�G,�E"�8ɓ���PPF��nJg�%G)���a��m�����ၕ�B���)L�5a�UyH�'�&����c6B��R�p�$�o�q�c9�����2ZFde�"{��E51�1M����<n�5h�~E�{P�j�y
ߓ5dy�3��l)
f/�	`�L� ��L�����쪡�N$��X�Idf��-O�<�(�%P�G[f��6�㍞�%�X�i*������_ ����0b��v3vn�#є��Z����Q�&����@dx����&DK#L�RT�KS�vAhiR̉�c#c7kvh!1��_�E��w$S�	ҳ�