BZh91AY&SYa}~ _�Px�׿�߰����Px�95 sFLL LFi�#ɀFM
{Jddi�      	D��O)�OS(�   ��y��sFLL LFi�#ɀF	"!�daLi�i4�hh  ɑ���@�RV�	��x�GաCGWbP
֒�aQ�V������I�?Rb���2�B�ŷCc;��!q���X�c'�`�
�dI8����
���NV����9�%�D�S��#s��1�:�����M�ax��D.�_�e�b�u�1♰˫���ʸ�Ɲ�m���6#Z�m��Ȳ���`ͼ�$�j�������@�D,Z25'�,�%$G�$�H\�l���i��Cj�I{u�ˏ�8���	H}r�ń����X�!HZ�]�t$<���o��^s1y�G*�yö���i�<�^A��öOI��������3�H*b�_�:$�h��t<l¶(�|#TFH�x�T�-P6��%��݆yxi("g�u�	�6T��(L��V��
Ｆ�X&�"X���S1f�T���܊�C\��ԇ aGam�	��% 'H�\�9Z���X,u�H�ȉ�Z騅4��c��a.�˂Le��i�(��O��H����0�����9��i��[y71�5ިE����&�E�D&�F̸P���9�A�Š.�p���a�Ty�6��ytcY��k&�H-�1���@o��� ����"F H V���d��m.�Zц욺��3��0yO<�S�����;-T*Xjb^
�;�G�mN��Ò٘�.��Gm2W�(����A�3 �"�Q�rE8P�a}~