BZh91AY&SY���u �߀Ryg����������`
�W�x�ף�4�㾾A��l�Q��J���Q�*i�OP��z����z��@�J�� @�M  �i&����i�4�&��H4�LL�0��RS�S�A��A�   4 JM��ة�(�G��G�#@�hA��� BI��&e	�L d 4 14:�UH���lX4�tUeU,�gK�Ѷ	$"L�� s���׮���;�a��R��5T��eTH^��luHTR���'4$��*!)��
T��K��ƫ��n@(�oDD6�u>�:�*��x��Ob�r��33bU�3ٕ�z�3�e�-���)c!�˘�Y��;�LQ����!�E�̉��&"$���#$�J�]c�Kc�eUR\c�ˬ��B�� �n�>�>G�U]��O:�m��GgR�y��Tӎǰ�����j�2�A�%�ƨ��6�� �����GҨ�
�O+��9嶻������Nc��%��{��� �0�����w\t�|O\a
�$�@�n&	��Je��C���=iO�TH]8ypOIX6����Ì4�D�ۜ"~����|s�����6fbd�E"M$�42��������B�xi91	d\Jܙ$�d!b�*s4�1w:4��rT0 %�m��҈�kuQ3Fd�2I(���;�擑��'�̱	'0�z�1�I7Վ�	2�T�R�ݱ��ڪ��̓�|��4�82nR�"�3$�%�M"xtm�,�H�" @���9�׬�33[�e�T����U�9v�X]�̌�"�eM�p�J.�W�#����	$�nߎB�F��i�l��qLF]�H��s}�V�w]y�̔@JR��C0��H�@L0J��1�:����Ӧ��u�f���I$�Ip�NŅ�''Ĺ�E�HHZ��2�M�՛�zR���	`�芆��y��'-�,�K��U�w!|	�r��#�0�UD�Y�g	{�7
l<�D��8M6-UU	C�?�s�n�\!
�$�I��ro*�Zz!F��LU�2�PaE@���Pp�b�*�ֵ�!��/1��!�ͳ�Lݬ�0�V���/5q-�����d��0�I&��j%@Z����۠�ͥd�_���<O���ʉ$�$5[\N7���k_������S6�a�JŕD�G(�r�ܫ4B�D�/�@�4Y3ԱW�bR�
 	+H�E/b-�N�/�S��P؆6��b��C���	##�*.î[�L�o�J[R�d���1Ŕ�n{b�L�E�N�r_=�ͅ�2n���1f˿����<!���r�VRKӐ�)�;�0l���x��)�T�1�Tk ��=� ���$�sYOl )6����jW/�TH59���OI��ǮWw�h�bFT�-Gͻ� fe��³}� (D`Lb(<�l��tD@�w�u���������_�6�Y�����lLR׃\�\�R�L��jR�&��IZie%�s�`��lO8��\˧����w��̥ʨ�+��3�����]L�����V抇������;0�9���cӴlu�6��*�oPS�6_���>�����>�����;n=BM�S�����OXi��'��}���i����f��M*�c�D)x�'��'CY%k_ {_-�qs�"�O�TN'p��;���'
C 6�D����"�Q�6ډ"�t���FU�ЮڗR�Ac�����\���P��TS�Q�0���>��s���?&���#�eQ!Q=���I�}H��Wt���$u�X�;{P���n��n�,��;��0� �1녌�0e t�<���'�t��Fz�:�*�k��U ��)�O	��t���Fl1+����*�TWw#�9��k�C����fz;;�{�QMr.��
�y��9����2�J.��B�=�ܖ0|�k�|�����C��%O[�=,��F@�ˢl�
�S����0DX[��3�
�` ���k,�Zd H�g/T�:�$"D[�8u*(�%�Y�[i�{8�R%��k�!n%���]��BB����