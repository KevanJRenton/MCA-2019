BZh91AY&SY��� �߀Ryg����������P>�wwt���[J�$�)��h&�SѤyO)�G�h=@y@�4L!&d@    �h��'���=G�Ch�b�M d�dɣ��i�0LM4��$MOCTأ�FT�j4ީ�2h  4yG���&�α\~�P��	+�S����9�>�@�F��m��۪����K\�8(dE��a�{)��i(�I5JV���uB(��bp�G��Z����˧�$���A��~�#��;�R
��9����U.�ǃ�(A��.��Jd�P�,���2����Lc�(+h��J�:ӗK�#��K�2�+d�JXٓ�Ν m�.��$nd�P���6�g�B��&�&Ȃ�/&�d�ܭ���U�"���ӍQ���HKKs�}��$D��)����j����[4fD���$�$���x�Ӕ��61?� ,E%4�!���"]�N�Zɐ�BPU_7Y%]D񚹥c��&����7v0��(2����469���}q�}GA�q�"w�����z!FZX'��e��p�C��HX�hR@�XY{�(J�*
���ivqf=��өLˠ�I�P2�����Z�="[G	9'��諺]\ä�8�m%���Ͳ1:�l�3���|�ٹw�*��S�{g���Μ1P��h�M��|&d)=>X��a�fwfsR�{�ݵ����ѺD��uhἲ�e�ӑ*()�Z)��Q

�E�2&r4��;1����c�<F!�&Ml)��2�ԡB��༤<�3u��]�(R�R���8��@o����m!	�}6_�d�If�� ύ�e�p��;�3&$`-�*]�5�������zeI��Hx��a�mH<�'�� gv��8�[a�L�B��#Ñqe	�tB;�S�@�L�LԔ���!<���\�Uk�t����0��I�C!'�h�-������p��h���4�7���4��&�;7O;�>����$�LG��Du�C,���"�5V'J`���ZZ9"Vl{��h�.�]��r�`��i�D����*��`�k@y���SCM(	&z��v{���=�qꥒ��j7����D��O' J��Yx�Q�����b�'tFy�����Q���02��\02�ƭ���֓E��5�Y�H,s��8��t���{����H~�ӎ%H�ab}S���2d���S2)SM;f����ڲJ	��d��څ���)���_P