BZh91AY&SY��$  �_�Pxc����߰����@ڀ�zOP12h    �����~��К4�  &�c�0L@0	�h�h`ba$"h���MM�A@��h�2f����E�e�$�2�1�d{�C�8�����Sb��0W��ُ�����cqb�2�R^zٛL��Yɸ�TŃ)�tG4Qb�$U{�W�5R��:o���3�t�ź��y���00�v�xw�&dnw71ӓуqi�3g!�)[mE:��_��7k�K$��$@�h^Au?�?v�(dX���
��s���Hp��!Fi�mJH����RE�xcz?C���ϨV-g.U��q�V�(��P�u���*al�p��d=�c㦚9����H�g����H�+39P[�x���|6CĄ~m�I���1S��I0,Fh��.���=�����$�%-u*��p�����ν�Bvۺ@Df�i��3��z�(���Ɔ�^0���N{u&�5J��!a�6
�?܈�E��Je��ur��:��ĕI�lŧv�[Q�s.1^�=�Yf��42���o]�gsc�p},���w!��u���γ�*"�Eb0@�2g[��e�>� _�ǥ�V�8��H����L�=k=��I��\HA�j�z��9���J���&0�-[tc�u�����~W�p���4���g���P�9܉�9��g�l�׹e���R]�e����)�bY����ɮ©tO	Y���\+����ᅆN����s�ِ��!_��%�IM�rE8P���$