BZh91AY&SYZе� k_�Ryg����������`      2h�14�@��`�M4 a2dшbi���4�&&�h �dɣ��i�0LM4��8ɓF!���`��i�q�&�CL	��14�@*�B4&	��@@&�4&���$�CA�$�@��#z�?W�dod��י/��X=�/#���յ�*�C$�T�~2Fi�L_�-a1!&��Q/�Q��5��#	iL#t�s�S��Χ��gs����N�M�֜q�-�R�R��Un`�*U)����.��g��}�=�%��gLے��v)����L���?G$�͞Y3�c�,ׄ@���E�����py�j}��R#�%6�텴�3LĦܾ7���F�o]!�+ʒ��"e3����#֔L�ɝr�h�b�T�s4�yu<V4I�OYȻ�W�6¡��J��5�Ζ`�]�T�6��2i�]�Y���BfZ�IL�����hM,�2y�=0�xC:��F2�$��,��)�h�����a�)�g�h��L�	C�k�SOZ�٭�YN���CZ��n����&s�Q�^���M9�۟�&ǥw�tR=X,����_�����,��mS���^
v��<�4��(�Mci~;�����c����d`�Ws������;F��O��yd��פ6��GĆ�)B=�(�4~M��n׭���=nQe?H���JR����%Ў�.��R�#�fzW�O����It�֔��{	���(��x�o���d�]��[+�"�]u��߯P}�����܌ux��ahS�Wo[/2Y:�X���c�Y�.���TSu��Yg�ڏl�?}�q�D�`��`�������O��^�fcS���KR옼�uw�7p�*%�txa8�҅�8�~�G4��b�,��))I#D.9n�2���N�c��d�DK���i�������u��bo]�Бͼ��bX���d�:�Dz��<�Q\ʋ�m҈����]��T�׌���{f�>4�
#kG�m!�b18.RJI$��$I(�X�QQ	y_#���h��QFL�F',"l��b-,ٛ��J�S�����aqNlc	���*�>�i���h�֡�.q;�OO�Iۨ��zDx�n�A��JCc��Ń�|�ۚ�H���M�c{z����ډ�K�L:�N�!܇z����v��Y�x����pp���	G(�t%EB^�����QcK\D>'sb�1&�IN��cU�&x�e�������X��^#�TGm�v5���N|��!'��Tm�����Whou4��&�
Os�%�ZV��S���u���!��c��I�S��խ���|,��ps�����3�a�2�f�r|��t=�}+���7q�5��w$S�	�X@