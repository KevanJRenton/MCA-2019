BZh91AY&SYQ֌' r_�Rxg����������P����\��c-	S$zDOSi��4i�hi�  6�  J��b�Ri�j2A��    %4$i4G�dɊf��h�SaOP�a��!�	�4ѣ4ɑ� �H�)��S5<�S�Si16���h  �ѓ,RLɍB��0�@��BWP������'�d��YL��$5l4U��P-�z �T���t f�C�����	���U޲&ʎ_Gf^/�Y�y�f��W�H�R���S�{9�\ws�r�;m֖7J�?�����(yN_����An��.o�$�4 $��^�ǁ�����b�.�¦2$!mс����trp:���	LHs��-),�*[h�	3\�M�Ѳ��T�\��CI�Ӛ2�����N
Mk�~v�bw�	"�q$�$�2x���:ô8z=�5��Jh�:�j�h�Zp��� *�!qALh£"�hE�Zurhs\A�
�H�Khc�\����8�<#�N�`����Y��rBY^�}�#3P���~���6啒B�>���KЍ�U[-��~e%�%�{pJyNV.UG�m��I`ߡ�r|v��zCA�H7�ui;�Ӭ��c
�G��O[�q�5����lR�<y	���K�&���<*������C33�3����W�oN�8�sc�ܽ{m6+��J	56X1d�Q�A,��e�j��~��E٘ӓ%sf%#���#=�"1M�:7N�v�ʓT���Ѹ�1���"�G*$�+>���-!iE�R�/4��A6�A8��Tm�.,Ϧ�J���M�N������.��b��;I���`��´bZb�B��QhW$�)��}�wq>��gbn�.:������vB@��t��
�b�HM�8,3ц��c+P�hh�5�y���/tJ N�ԛL�/����U*�r����B)���+����6�w�I�$aa�F�sf�>0;����;@�Vg�.��vo$n"�h�B཭u�t!Z?���^#p�V̷�.�00bAT�p�cot�9�����Z5�B)Db`ɟ�3�Q
�mLj*^��?`כ֨\���A�qR�n��]"���D�d�M��]x2�_$����@hO,t�e*�{��?��t�"����ka��(��v�4h����1�R
X�d�1�snT�-Eـ��.�p� ��N