BZh91AY&SY'�W �_�Rxg����������P��[Ɉ��M4%
d&�M&��Sڞ�z��6���F�PPp�L�FL0	��bd4���	M
h��m'�d�4Ƃi�@   4�#��i�`��244D�&�i�iQ��S��)�� P����I6�s
��b�
`�����/�Ak�����>��s��0��d����(u��JL���W!*0$�_�r
�?��cFZ����Ͳ�G�R6���lyb/UB��[�w�T���<s��u��J69���p�M��VNE�<��P��^��{�H�A _2� -F�I�Cu���OةT��F���/;V`K@R��ٱS����ʃ��Bw�[	���1�!ph���ٌ���B��s��z�)-C2r̙E4
Z]�����6���ƃ�n$�ē���a<	�rn����_�AEP���"
�H�w�KBd;�A�ҧ�ӄ�L՝f@\�v1M�t/n�Kan�`��^���_������ק�P�u2L�ol����>^�/���,b��gE�QM�:9*:�U"�=5p~F~=O��&ϖ�W�e�bJ� �Mj�G�!`ʊf�HB��Z:/�%˸6�]��A�i���|�d��OZ<c��O�J��4i^�R<="i�x�]8�&����2�u���C33�3���,���0R��	�]���ګޘh�;�U���R�*yd�����C�S�и��uW���\4s2)��QN�B3�o�f3�'��󔮾�h�&y��xjV�5��9Ad���k261�tL�uaH�p�i�5�l��j(i"��kȝ�85pO1$���F��F�ͭ:����wV���TA������N�2ÍK'hXZq�K�r3e ���@��p�i������n O��N5������uF����a'm���BP:e���J+����r��w��S��,,e-��3�{N����:�r�&��ZR�k�U@��۱y�9��q�H�K/4�V�L�؆7b�\�d5���j���XM��xF�K=�  ���M4�$���@�i��$f. ��D�b�����ک"�޽�aS`�徏K�%���d��|�hӜ����\��.d��fF�h6['�%�����U�����Gg���1���0%�v{3�hD�KRh΃]�Jo��#�:�U�S�e�qZ���ip'������)��=R�