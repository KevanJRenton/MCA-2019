BZh91AY&SY��s _�Rxg����������P޸�c��w9Ҵ�ДHĦъm hѧ�i�@��4��*~�ئj41      %4"A�L��F#M�d4 ��4��a4�C �a&&CL� �!)�&�S�OI�z����F� !��I3&5�gф�D�1��D?|�	�c��f�˝�>}����~�YC�Qe V��5�3Q�w�5��[�(�gADB�`�6wxqr?ֻ8��̓g��0T�?��u?#�ja�q�͑���ӡ-ۨ��u*S V����&n@��=�I�H +�8	#�a��<�0��1c�+lFfa�mzq9��ua�,�'&����7��s���F2\L,J�vc�p4��)��	F%TQy���h�U��~��m��<FD�{��t�\��@�j��8C�9Mb
�	)���a�[P]�HDv\H8"�Fڋ��CT��a}�jm��m�;%}�+����bW��+U[%R�<^�j
=����(�'�;�t0�B�v�ެ�0b�f0	�Ӏ��Ed5.�m�$�o�dp_�42��:��!�uCT!0%KS~Ht@16S�� g�26T�Q�CT����zui�����q��{��Hpu1�aY�J�t�M>0$�A�t�D�m��4<�&�C33�3���1n�n.]���BhX�鳁a�1�9AhWC i��N�K�����%���������eҊ�:r��	���F��<��rW���hQ�}6�Lhe|$�p��[V�2~˺H\(�l�V�A���Ą�����Kn/�dU�"��7��/5#���t���Q�,�Lk����=h+�s�3f��D�gu3��|]��&*��:�gp�E�Ұ���V��y�"f���H���L�((����$,tbjT2��u���0JH�;�}6���2lZW5ri���(�d�#dU��Ĵ��8�d�E�2<�"�:	��T��c�X��$��h��p/�tm����²�ֺع��?�9��1�T��@_ 0``�AV�p�c���Y�ע�c6}[��VF0L�N��2Q��EZ����VjA����[�%���i*�R6fщ`��&eA� QS�����{h-z�p��u��T�v�x����Hx�i�d�D� �TI% a/[kJ�2��F�9Yt=��&�F�#2Z��o���)����