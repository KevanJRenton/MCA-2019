BZh91AY&SY���� ߀Px����߰����P~t.l@G4d���`F�b0L�`�4�H�dzS2LCFChP(
i�驦�SC� �  �sFLL LFi�#ɀF	MM4	<�Sl���C�Tf�(�J�!!��cRhm�B��w��~�"��ah���rΨ���὜ķ-k�RY��&s%ժ�iC���������9���#TJ� `M���e����z��1KuJ��+�c!����.&ͭY���ơ5�dQ�fA~b7��'�/��,�Ɯ��dr�9�����p"١�fہ�&F�����(!�EfK
U ����ȃ�UF!J�(9C�lfh����=w�Bƶd��7���$(R��{��~9�)�#�����!,V�!嗩y�͞�AS��t�zC���_�҃Q!�	�s�&�f�?�U�R| ���fz��E�A�T�M���I���*!\�.]��A�A�t-��Z0��˭��|h�
�%�V�@}wS2><��/q���؟0�az�KH�l��-��%܌��������;l��Z�zIL 
���Uh]n���َ����>� ��%lΌ�Չ��KKB��$��QmB4·E�"�X"��� [�[W:���t����J�dj�E���&%��R�Q��4f���v �ZCW:���C�.>��;@���"�v�{�J���ڎ>�� 8����	H>���;vԩ�
��"�"X���A�{$!)�dS�a���)�#��3D��P�)���d]a�$DV�ׂ?��B���#�*y����y��d���lV�s)�z6�p�����.�p�!ї�8