BZh91AY&SY\: ߀Ryg����������`�  �   dɣ��i�0LM4��8ɓF!���`��i�F��oT4�@� �d@� 8ɓF!���`��i�q�&�CL	��14�@H� �4 SA2M=F�ڌ�m��$�0t��?1��1WKY4/�CĐ��	���������~I��.,s�#VV�2B���'{A �?�1���X��@H,	�F�|�^����Q4�G�hť�K����4����\J݂�[�ȢpR�"�B���a)��MZ~bL��:/�A#�E�B'K{��mƮP����%5�2x�Y2��j �T��8+�|iݳ���T4�|=A�I�U�Nd�:� lʊ����>ԸX4�{~f�_�4`�{sG>)�L|x�?�\נ������傳'��AF����î�����Л�`�r4ha�}�n���[�r���]�pt�CM�L�e}L�6��C�؉�����}h�+#�t)���3�ly�m��cp�M��~`q��Gh�����X����̨4�2�[�������(�2X�H�~��f�K�	�"�y,dCL,�I
�b���Y�`�l����$�Nɫ����Cp��Ͷ�p	 ��lZ���į��Fr"�e0
'0�	P�0��*bO����N���N]_2�P���]ӆ���]�/��Fb�.�\o$�!�SW7yP�SY�S!Sq3���X��_.�2���8J�@1�=~'ƀ�!�l l?DB$�?|�֓��i<�݀�Z�#��G$��Zϵ��B��}~��$[A{��'��#QY�?n#�V��t�"��z/G�=����)�M$h+�w��L�U��D|<et�H �2d�	Ϧ��P�����y��,�H�b�_�WS.Ε#�e�	�D�&��;��QT�J�A41)�!UaMB��k����;0*�.DQ[�`q��� �F�������pF͡e3�HkG�J�B�_�ė�̂��}X��)�*z��騧��
���pKA.TP�GT�"1$1�4��z?�9�cF�
�>�p�4��ML��rK��>���+�7���qD�����	4%����ʪX61z���[D�U�O�.$"�x�b�J�7�孤�����$�϶̙�:+λĥ��_S^��čb����qP*-��j�g�1���@�:ks[K	,�(5P�~� 9�Ɂ'��h!1I�'
5ʘ��T,�E�Ћ�&� .CAL�J �.�W0�
P#)�g_ ��@�΄�N���(@��j@�u�S/���C�/b��fdi5����`yl>&�LH�Ѱ�5k��2ߏ2\��@`{D/A����*{�a#�v����5��a��6-�#́��s��� I^K���gE��`�&��H��t�Az(Y"Ʌ�hs"GR��%TI�{N�3K�� ����R*`��p�.������M�ix��o���4�&�J����:�5��^lJ�35�]W�\L�`+�Ӭ��әp#Y��fi0<O�a4��D�B�F$K���@ja�(�̈[p���޷��+4а�)"�a���}vx���6��0�ױ ���H�
��@