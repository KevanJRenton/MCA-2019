BZh91AY&SY�OO� �_�Ryg����������P������U�Q&���Q�i �� ���J�'����4�&��M4�L!��4 �C  �Є&�����e=A��j4  �2dшbi���4�&&�h �	"	�LSh�S��Sjm�SLh22�0�I�o��A%D��(�y8c4�}S���phe�p��@GE�H��(F��D.(���@C�@�ns��3�z�8b��.�6?ֱ���u!6�H�����x����)�wslm�;j�Y�#X�AxE��D�`��tWk�Bc%Bi8�F FB. ec����!O.�Կ�4e�=iX�0���<�x�%�����a���$���M�f6�I���Z��/B�t����o�`�ŝ�-����R��>5ʩ{nsX�*p�8L���#q$�$�l'�9^��������5U%4� ���w㝈�L�zq�^E jfzb��6������*��Ί�\Fl��3J:��������)�X�UwLO=Oe{�ݗhU��͊�%��6���9T��.��7��I�f���.���;fw�m*%�$L��#�{@�D���Bt�;�����A��]� ���X|��UY)�R��m(X�5��U���-ʙ�4�}���4��8OVk�42��lZP�����t��z���2�rpD&ߐ�ՏWM��v��(�){՘��� �wg�d<GbL�%tQ/�d�h�R5��"]�t\����W����MqO�˸�R!��2Ҭpd��k�2i��s�g9��esć���@d�AN"��%ӓ����T���#	�Q�{�^3�T����gdƼ�պʤ�Z�����Q��v��*�C�a�&8L5�(m�Q.�.#��)`2�<4
���d��2&��iM���Τ�3���϶f��bP�0E���� ��ld�f�9���4�94�w��00��F%d,��N���Z�i���ЙM�*��M����y��`.b��IE �܏0X��I�ucb�X�:�Y���L=e�lsΘ����2`�<b�2NQ���cj7� V\%�|�P�ҘŠ��c����*a�Zw,)���]Sΰ�Q���w��h�[�)�e�%,�+.�����F´kb��;o¨cY ��vSA���G���1���0���6�^�LT/��Y�N�ّb���,�X��g�Dv�fKy�!�rE8P��OO�