BZh91AY&SYw�<�  �߀Px����߰����@m�
Jz��&�L&�L�24 �0�=L��h@@i��sFLL LFi�#ɀF	M4#F�&��M�z�e2 ���&���]P�B SH�P���=�_�&��=�D0��H�4.�M�l�]����y�����ɕЁ�t������T�+��q[-f�G�XBI� ��l��m����OOgi`�=������3����m�d�Y蒥�|�V���:�Ta�5{��{���J��28�3{�b-�g��#�L�������H�jt�L�D�B�
4�f�"���8��9Ӛ�!
��;�G�V�Q���ҦR���ai��i�k���cm(ӡ& �v��Y��B�h���d@�b(��Y�]���bύ��c�8��s?!wx�:������X�T)0͕��@3V�~}�$ئ����\RC�y����9��Jʼ�+]Z�Fuנb��
�߱?��U�����(z�
�̗j4^��\!s��r	��/�Hz�MB.��g�z�Zj^T�,M�0���G���*�tfXf8O[H�s]��V������%��Z#Q�"54�v@;���*>��r�dR�V6@�Ɋh��W\�Q%�BR�,]�:M'���$�}�Pk��׭����~&���M���z�g���A�7#����.cb���H��W��wZZb+BET������yoF8���� .J��OT��IZ�'@�=���ԅĊE,4���AmEb#���G�)����6Ѱ��e?wx�����_�.�p� �y�