BZh91AY&SY��.2 �߀Ryg����������`�  
     ����F��f�1h � �8ɓC�� �� �M4i���&MF&�04ѦF�c��41�0�L �F��2d��bh�#0�0Mdh$M4h&�i���j�� z�1���SU�L ��0P�	��H>qFe|���&�a4"ۏ��#����2����O�,m�d�y�P,]�M#��#@Ԙ��
ā*0	 ūA2IXhg�B�h�<�
&�b�ɥ����2���̸��Ѵ����T��mH%�R��Ozj��I�Y�B��( �z�_�h[��DAtY��%�%= lpe'���*8�y�9��۾2ݳ���T2��z�H����'2a�� 4�a0r�ؗ!������óo�f������#LL|y���h-W�rK��#.<�V3�MɁ0(��ŻR�u[�xA���`6�47�#�ﳀ�O��K໠u���!��jʴR	�$I���!��Dԕ��{�UT�Ǜj����8����r�"n�m�ߜ�@\w��=����H�BJ̨4�2�[������&U�-M>�ߌ��0�)��"�Y�$�4=�(b@`X����	%�vM\0	��n�f�nG @�0 X����_o�kd��`� `�o�D�B� ?9B@n�#��)*���e@����]Ն��d��/5��4(�.{����6�j��*�h5�
�EC��$�Z�W
H�.��gu���(jV�pcj{<V�@Y�;������0�u�ڵ)-G�[��yA�ʤr�5����R2X}_^ �����}�2+2G��ƟJ̼]�������K�SHMį3���S>��p� Ƞ\�b&L�>�s�p�@]���<�4X�"I�I9uSO_J�@˱&HR(��)Т�E()�Ц( �U�Y5
K�ז�%����K,�2*�>���BJ̍�UQˈ:�E�w��6a�<��'�4X��I�V6�j=��.��Q}e�.���zb9�@��G�(��#CcL�\Wx}���4j �IAϑ�4��M(5#�p�i�|Sq�+�3C9�%�7���$H�.!��}<���a3@��]�R�&��)>и�=%��@��p�@nNc��$@��׊�!2�Q�Iɨ��`b`
ZnB���^������� x���N���}�`��H$#�@&�hֶ��@���c�P��~L	<Ri�$�@@��&(�*Ӧ�\<BĮI���D>%\^+��S(���>��@�� ��Jx��c����$�)��4CRc@e�8)�P��޶���#�k��-F���6�@��v��r�����.��R  (�����*~CXH�<��=��k3Xg�҉ �����LD$1{�u��p^sa5 � �AyT� ��rarL_F�S&�@hd��5�:��e��7G�MH��S����%e�6�ю�hn�*$�q�W3@L3�k�cX�;�͂�ƍF��5׆��f�@�KVd���$dm�&�����TH[�p�� ��щ�A�5�F��<&�l7��b���4,$�H�Xq0_�m�cVᔘǔ$�%�%�؄b����)��q�