BZh91AY&SY�ӧ! �߀Ryg����������`  
     �(�M b   � ��4b�` `M0F	��� 0�2h�14�@��`�M4 a2dшbi���4�&&�h �dɣ��i�0LM4��$hL�2d'�2&CG�Ɇ����	&�:AZ�`�$%jBZɂ����<���w܄I~��M���S���S����jՍ��HW%�����?&�`5&)�B��%F �$BU�����[AD��b=�F,�^~>��<�'3�-%gb9�=|N��),�l��T�?Ț�~d��P�t
!R.���gO���6�G(g`vJ�Md�3)<�,�Q����o-4(Wo%�����:�t�}I��\��L5U fTW� [���%����2�3�}X/�0v��#,1bc�m�����-Io�`���u�Ḿ0(�������PU�^Paz	is�a��H���J������-9�Β8��!��������D����LqGx椭N��P�u�~�#w�Chz@�٨��6�m���C -=\�Ob�m�$|BH���&Qˑ�Ark�\�
*̖M?S�3���Eİ�L,aI"�b���ƕ��m�ir��W�bjрMۋp��F�r7� ھ�����%u�"�3��`�0+ �0�|��"1L0#G#��� ��*
B�;�a�7�+gUڪ���;�W����@��$��!�S_IP�)���S1Sq3~J�/�����U����;�����m`zO꠿��-6�@
H�j��$�<��x�PG�pR8H��|�vA
Fj���E�	�����gL��#2�$ɍ�-��\�'���r=��qj�XW0��[ ��\)��Ҭ!@2��z�l�A2d���E}�o��;ֈ,X�"I�I}��]}*K�e��$(��$S�EP�P$R	��LPA
���5
KQ5ۮ�E���Kk�(����0�!%VFҪ��:�E�6��g�Xmj@�6����!Xz,m�S*T����QO�v�*���#�,H�p@��H�y!�1�uSp~����4j �P����R%4,�ԏD��8��x�Ӑ���b�����Z�	3K�mZ�F�������h-��m_��Iȴ^(�.��s�Ĉ����W�	����N!�W��,a�.���&�+�� ���N���|�`��H$#�@&��Z�X	i�U
��Qn�)`~L	;����p� C\�\K Y�r.Aa+�j�4ϰ�Bۅik
`�/�l:�W���{�*p��P�$ULԁ��3Lh��|�>b��n�Ff�`ř�m��k0��5ky]h9V��R�jD�������§� �$}'`{2F���4��Ŵ�H;�b`���� I^K�����;	����t�ApyԵ"��Ԙ}�H�T 0d��5�q�6�Zu�9�=��EL r�.��4q(�,�nZ��7���gD�n5*�`(�t�kS���+��h�aluݡi3ax�	���b�V���5���?��e�*
$-��`�o �;���A�5�FEV��l9"���X�B�L��U�W��ϖ��Vᔘ��_a0cIt���FK���"�(Hk�Ӑ�